`include "defs.vh"
`include "timescale.vh"

module core_pipeline(
    input rstn,
    input clk
);






endmodule
